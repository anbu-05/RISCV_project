module sram_tb;
    
endmodule