// module RISCV_core(
//     input reg enable, reset, clk);

    