module top_tb;
    